/escnfs/courses/fa22-cse-40462.01/dropbox/cgillila/VLSI/muddlib.lef